* Simple NMOS Transistor Characterization

* Include the IHP PDK MOS library
.include /opt/pdks/sg13g2/libs.tech/ngspice/models/sg13g2_moslv_mod.lib

* NMOS Transistor
M1 D G S B sg13g2_lv_nmos_psp L=0.18u W=1u

* Voltage Sources
VDS D 0 1.8V
VGS G 0 DC 0.9V
VBS B 0 0V

* DC Sweep for Id vs Vgs
.dc VGS 0 1.8 0.01
.print dc I(VDS)

* Save all results to a .raw file
.control
run
wrdata output.raw all
quit
.endc

.end
