* Device Characterization
.include "/opt/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib" mos_tt

* Supply and Biasing
VDD Vdd 0 1.2
VGS Gate 0 DC 0.5
VDS Drain 0 DC 0.3

* NMOS Transistor
M1 Drain Gate 0 0 NMOS L=500n W=30u

* DC Sweep VGS
.DC VGS 0 1.2 0.01
.PLOT DC ID(M1)

* DC Sweep VDS
.DC VDS 0 1.2 0.01
.PLOT DC ID(M1)

* Operating Point Analysis
.OP
.END
