** Simple NPN Transistor Amplifier

.option TEMP=75
.option warn=1

* Define power supply
VCC Vcc 0 DC 12V
VBB Vbb 0 DC 1.5V

* Define the transistors
Q1 C B E 0 npn

* Define resistors
RB B Vbb 10k
RC Vcc C 1k
RE E 0 500

* Load capacitance
CL C 0 10p

* Define input voltage
Vin IN 0 SIN(0 1m 1k)

* Coupling capacitor
Cin IN B 10u

* Simulation commands
.control
tran 0.1us 10ms
plot v(C) v(E)
save all
write $(RAW_FILE)
.endc

* Include standard NPN transistor model
.model npn NPN(IS=1E-14 BF=100 VAF=50 RC=1 RB=10)

.end
